/***************************************************
Student Name: Yu_Ho_Chang
Student ID: 0716046 
***************************************************/

`timescale 1ns/1ps

module MUX_2to1(
	input  [31:0] data0_i,       
	input  [31:0] data1_i,
	input         select_i,
	output reg [31:0] data_o
    );			   

/* Write your code HERE */
	always@(*)begin
				case(select_i)
					1'b0 :
						data_o<=data0_i;
					1'b1 :
						data_o<=data1_i;	
					default :
						data_o<=data_o;
				endcase
	end					
endmodule     
          